// -----------------------------------------------------------------------------
// Universidade Federal do Recôncavo da Bahia
// -----------------------------------------------------------------------------
// Author : João Carlos Bittencourt
// File   : selfcheckDriverVGA.sv
// Editor : Visual Studio Code, tab size (3)
// -----------------------------------------------------------------------------
// Module Purpose:
//      Módulo de auto-verificacao para o VGADriver640x480
// -----------------------------------------------------------------------------
`timescale 1ns / 1ps
module selfcheckDriverVGA();
   logic hsync, vsync;
   logic [3:0] red, green, blue;
   initial begin
      fork
         #00000 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #00030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #00070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #00110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #00150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #00190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #00230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #00270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #00310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #00350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #00390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #00430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #00470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #00510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #00550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #00590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #00630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #00670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #00710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #00750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #00790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #00830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #00870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #00910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #00950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #00990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #01030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #01070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #01110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #01150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #01190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #01230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #01270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #01310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #01350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #01390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #01430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #01470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #01510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #01550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #01590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #01630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #01670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #01710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #01750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #01790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #01830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #01870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #01910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #01950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #01990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #02030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #02070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #02110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #02150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #02190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #02230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #02270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #02310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #02350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #02390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #02430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #02470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #02510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #02550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #02590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #02630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #02670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #02710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #02750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #02790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #02830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #02870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #02910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #02950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #02990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #03030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #03070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #03110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #03150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #03190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #03230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #03270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #03310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #03350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #03390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #03430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #03470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #03510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #03550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #03590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #03630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #03670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #03710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #03750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #03790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #03830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #03870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #03910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #03950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #03990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #04030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #04070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #04110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #04150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #04190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #04230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #04270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #04310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #04350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #04390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #04430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #04470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #04510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #04550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #04590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #04630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #04670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #04710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #04750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #04790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #04830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #04870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #04910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #04950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #04990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #05030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #05070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #05110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #05150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #05190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #05230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #05270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #05310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #05350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #05390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #05430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #05470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #05510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #05550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #05590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #05630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #05670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #05710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #05750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #05790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #05830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #05870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #05910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #05950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #05990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #06030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #06070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #06110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #06150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #06190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #06230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #06270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #06310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #06350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #06390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #06430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #06470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #06510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #06550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #06590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #06630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #06670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #06710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #06750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #06790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #06830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #06870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #06910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #06950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #06990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #07030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #07070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #07110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #07150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #07190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #07230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #07270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #07310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #07350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #07390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #07430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #07470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #07510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #07550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #07590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #07630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #07670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #07710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #07750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #07790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #07830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #07870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #07910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #07950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #07990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #08030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #08070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #08110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #08150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #08190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #08230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #08270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #08310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #08350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #08390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #08430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #08470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #08510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #08550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #08590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #08630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #08670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #08710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #08750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #08790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #08830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #08870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #08910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #08950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #08990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #09030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #09070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #09110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #09150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #09190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #09230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #09270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #09310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #09350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #09390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #09430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #09470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #09510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #09550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #09590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #09630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #09670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #09710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #09750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #09790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #09830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #09870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #09910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #09950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #09990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #10030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #10070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #10110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #10150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #10190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #10230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #10270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #10310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #10350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #10390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #10430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #10470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #10510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #10550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #10590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #10630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #10670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #10710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #10750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #10790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #10830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #10870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #10910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #10950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #10990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #11030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #11070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #11110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #11150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #11190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #11230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #11270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #11310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #11350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #11390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #11430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #11470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #11510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #11550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #11590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #11630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #11670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #11710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #11750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #11790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #11830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #11870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #11910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #11950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #11990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #12030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #12070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #12110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #12150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #12190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #12230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #12270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #12310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #12350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #12390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #12430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #12470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #12510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #12550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #12590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #12630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #12670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #12710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #12750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #12790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #12830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #12870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #12910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #12950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #12990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #13030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #13070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #13110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #13150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #13190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #13230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #13270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #13310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #13350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #13390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #13430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #13470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #13510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #13550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #13590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #13630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #13670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #13710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #13750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #13790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #13830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #13870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #13910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #13950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #13990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #14030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #14070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #14110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #14150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #14190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #14230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #14270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #14310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #14350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #14390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #14430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #14470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #14510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #14550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #14590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #14630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #14670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #14710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #14750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #14790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #14830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #14870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #14910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #14950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #14990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #15030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #15070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #15110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #15150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #15190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #15230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #15270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #15310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #15350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #15390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #15430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #15470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #15510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #15550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #15590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #15630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #15670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #15710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #15750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #15790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #15830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #15870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #15910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #15950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #15990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #17030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #17070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #17110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #17150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #17190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #17230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #17270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #17310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #17350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #17390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #17430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #17470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #17510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #17550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #17590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #17630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #17670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #17710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #17750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #17790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #17830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #17870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #17910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #17950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #17990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #18030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #18070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #18110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #18150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #18190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #18230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #18270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #18310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #18350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #18390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #18430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #18470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #18510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #18550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #18590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #18630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #18670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #18710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #18750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #18790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #18830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #18870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #18910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #18950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #18990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #19030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #19070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #19110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #19150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #19190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #19230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #19270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #19310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #19350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #19390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #19430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #19470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #19510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #19550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #19590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #19630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #19670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #19710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #19750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #19790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #19830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #19870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #19910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #19950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #19990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #20030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #20070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #20110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #20150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #20190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #20230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #20270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #20310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #20350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #20390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #20430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #20470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #20510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #20550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #20590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #20630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #20670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #20710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #20750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #20790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #20830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #20870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #20910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #20950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #20990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #21030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #21070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #21110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #21150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #21190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #21230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #21270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #21310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #21350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #21390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #21430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #21470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #21510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #21550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #21590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #21630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #21670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #21710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #21750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #21790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #21830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #21870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #21910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #21950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #21990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #22030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #22070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #22110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #22150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #22190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #22230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #22270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #22310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #22350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #22390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #22430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #22470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #22510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #22550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #22590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #22630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #22670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #22710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #22750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #22790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #22830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #22870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #22910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #22950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #22990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #23030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #23070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #23110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #23150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #23190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #23230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #23270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #23310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #23350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #23390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #23430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #23470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #23510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #23550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #23590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #23630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #23670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #23710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #23750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #23790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #23830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #23870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #23910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #23950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #23990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #24030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #24070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #24110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #24150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #24190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #24230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #24270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #24310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #24350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #24390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #24430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #24470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #24510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #24550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #24590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #24630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #24670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #24710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #24750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #24790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #24830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #24870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #24910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #24950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #24990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #25030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #25070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #25110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #25150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #25190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #25230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #25270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #25310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #25350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #25390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #25430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #25470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #25510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #25550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #25590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #26230 {hsync, vsync, red, green, blue} <= {2'b01, 4'd 0, 4'd 0, 4'd 0};
         #30070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #31990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #32030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #32070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #32110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #32150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #32190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #32230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #32270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #32310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #32350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #32390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #32430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #32470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #32510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #32550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #32590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #32630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #32670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #32710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #32750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #32790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #32830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #32870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #32910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #32950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #32990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #33030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #33070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #33110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #33150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #33190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #33230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #33270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #33310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #33350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #33390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #33430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #33470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #33510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #33550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #33590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #33630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #33670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #33710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #33750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #33790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #33830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #33870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #33910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #33950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #33990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #34030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #34070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #34110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #34150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #34190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #34230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #34270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #34310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #34350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #34390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #34430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #34470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #34510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #34550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #34590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #34630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #34670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #34710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #34750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #34790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #34830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #34870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #34910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #34950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #34990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #35030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #35070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #35110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #35150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #35190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #35230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #35270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #35310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #35350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #35390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #35430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #35470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #35510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #35550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #35590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #35630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #35670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #35710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #35750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #35790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #35830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #35870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #35910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #35950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #35990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #36030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #36070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #36110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #36150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #36190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #36230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #36270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #36310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #36350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #36390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #36430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #36470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #36510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #36550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #36590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #36630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #36670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #36710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #36750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #36790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #36830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #36870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #36910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #36950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #36990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #37030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #37070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #37110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #37150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #37190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #37230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #37270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #37310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #37350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #37390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #37430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #37470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #37510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #37550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #37590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #37630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #37670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #37710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #37750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #37790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #37830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #37870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #37910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #37950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #37990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #38030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #38070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #38110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #38150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #38190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #38230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #38270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #38310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #38350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #38390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #38430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #38470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #38510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #38550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #38590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #38630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #38670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #38710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #38750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #38790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #38830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #38870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #38910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #38950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #38990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #39030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #39070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #39110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #39150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #39190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #39230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #39270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #39310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #39350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #39390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #39430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #39470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #39510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #39550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #39590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #39630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #39670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #39710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #39750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #39790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #39830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #39870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #39910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #39950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #39990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #40030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #40070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #40110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #40150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #40190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #40230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #40270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #40310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #40350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #40390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #40430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #40470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #40510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #40550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #40590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #40630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #40670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #40710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #40750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #40790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #40830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #40870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #40910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #40950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #40990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #41030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #41070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #41110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #41150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #41190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #41230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #41270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #41310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #41350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #41390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #41430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #41470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #41510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #41550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #41590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #41630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #41670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #41710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #41750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #41790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #41830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #41870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #41910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #41950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #41990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #42030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #42070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #42110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #42150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #42190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #42230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #42270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #42310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #42350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #42390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #42430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #42470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #42510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #42550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #42590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #42630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #42670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #42710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #42750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #42790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #42830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #42870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #42910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #42950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #42990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #43030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #43070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #43110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #43150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #43190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #43230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #43270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #43310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #43350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #43390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #43430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #43470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #43510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #43550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #43590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #43630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #43670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #43710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #43750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #43790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #43830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #43870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #43910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #43950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #43990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #44030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #44070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #44110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #44150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #44190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #44230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #44270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #44310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #44350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #44390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #44430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #44470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #44510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #44550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #44590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #44630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #44670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #44710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #44750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #44790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #44830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #44870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #44910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #44950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #44990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #45030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #45070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #45110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #45150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #45190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #45230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #45270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #45310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #45350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #45390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #45430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #45470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #45510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #45550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #45590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #45630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #45670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #45710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #45750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #45790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #45830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #45870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #45910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #45950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #45990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #46030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #46070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #46110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #46150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #46190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #46230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #46270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #46310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #46350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #46390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #46430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #46470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #46510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #46550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #46590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #46630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #46670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #46710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #46750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #46790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #46830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #46870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #46910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #46950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #46990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #47030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #47070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #47110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #47150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #47190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #47230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #47270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #47310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #47350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #47390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #47430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #47470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #47510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #47550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #47590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #47630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #47670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #47710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #47750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #47790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #47830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #47870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #47910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #47950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #47990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #48030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #48070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #48110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #48150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #48190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #48230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #48270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #48310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #48350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #48390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #48430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #48470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #48510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #48550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #48590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #48630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #48670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #48710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #48750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #48790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #48830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #48870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #48910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #48950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #48990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #49030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #49070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #49110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #49150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #49190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #49230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #49270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #49310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #49350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #49390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #49430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #49470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #49510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #49550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #49590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #49630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #49670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #49710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #49750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #49790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #49830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #49870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #49910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #49950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #49990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #50030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #50070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #50110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #50150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #50190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #50230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #50270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #50310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #50350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #50390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #50430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #50470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #50510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #50550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #50590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #50630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #50670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #50710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #50750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #50790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #50830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #50870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #50910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #50950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #50990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #51030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #51070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #51110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #51150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #51190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #51230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #51270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #51310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #51350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #51390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #51430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #51470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #51510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #51550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #51590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #51630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #51670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #51710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #51750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #51790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #51830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #51870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #51910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #51950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #51990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #52030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #52070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #52110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #52150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #52190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #52230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #52270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #52310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #52350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #52390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #52430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #52470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #52510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #52550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #52590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #52630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #52670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #52710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #52750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #52790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #52830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #52870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #52910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #52950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #52990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #53030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #53070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #53110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #53150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #53190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #53230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #53270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #53310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #53350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #53390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #53430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #53470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #53510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #53550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #53590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #53630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #53670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #53710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #53750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #53790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #53830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #53870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #53910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #53950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #53990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #54030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #54070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #54110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #54150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #54190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #54230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #54270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #54310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #54350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #54390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #54430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #54470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #54510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #54550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #54590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #54630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #54670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #54710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #54750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #54790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #54830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #54870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #54910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #54950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #54990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #55030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #55070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #55110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #55150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #55190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #55230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #55270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #55310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #55350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #55390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #55430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #55470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #55510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #55550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #55590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #55630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #55670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #55710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #55750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #55790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #55830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #55870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #55910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #55950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #55990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #56030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #56070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #56110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #56150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #56190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #56230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #56270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #56310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #56350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #56390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #56430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #56470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #56510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #56550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #56590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #56630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #56670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #56710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #56750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #56790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #56830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #56870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #56910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #56950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
         #56990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 1, 4'd 2};
         #57030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 5, 4'd 2};
         #57070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 5, 4'd 2};
         #57110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 9, 4'd 2};
         #57150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 9, 4'd 2};
         #57190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd13, 4'd 2};
         #57230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd13, 4'd 2};
         #57270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 1, 4'd 2};
         #57310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 1, 4'd 2};
         #57350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 5, 4'd 2};
         #57390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 5, 4'd 2};
         #57430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 9, 4'd 2};
         #57470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 9, 4'd 2};
         #57510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd13, 4'd 2};
         #57550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd13, 4'd 2};
         #57590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #58230 {hsync, vsync, red, green, blue} <= {2'b01, 4'd 0, 4'd 0, 4'd 0};
         #62070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #63990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #64030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #64070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #64110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #64150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #64190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #64230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #64270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #64310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #64350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #64390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #64430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #64470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #64510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #64550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #64590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #64630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #64670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #64710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #64750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #64790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #64830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #64870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #64910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #64950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #64990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #65030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #65070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #65110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #65150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #65190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #65230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #65270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #65310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #65350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #65390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #65430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #65470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #65510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #65550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #65590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #65630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #65670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #65710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #65750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #65790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #65830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #65870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #65910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #65950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #65990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #66030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #66070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #66110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #66150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #66190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #66230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #66270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #66310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #66350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #66390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #66430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #66470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #66510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #66550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #66590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #66630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #66670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #66710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #66750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #66790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #66830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #66870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #66910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #66950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #66990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #67030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #67070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #67110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #67150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #67190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #67230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #67270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #67310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #67350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #67390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #67430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #67470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #67510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #67550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #67590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #67630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #67670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #67710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #67750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #67790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #67830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #67870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #67910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #67950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #67990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #68030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #68070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #68110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #68150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #68190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #68230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #68270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #68310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #68350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #68390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #68430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #68470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #68510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #68550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #68590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #68630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #68670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #68710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #68750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #68790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #68830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #68870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #68910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #68950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #68990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #69030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #69070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #69110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #69150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #69190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #69230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #69270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #69310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #69350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #69390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #69430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #69470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #69510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #69550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #69590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #69630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #69670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #69710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #69750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #69790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #69830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #69870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #69910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #69950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #69990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #70030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #70070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #70110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #70150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #70190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #70230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #70270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #70310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #70350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #70390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #70430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #70470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #70510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #70550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #70590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #70630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #70670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #70710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #70750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #70790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #70830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #70870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #70910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #70950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #70990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #71030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #71070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #71110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #71150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #71190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #71230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #71270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #71310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #71350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #71390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #71430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #71470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #71510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #71550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #71590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #71630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #71670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #71710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #71750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #71790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #71830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #71870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #71910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #71950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #71990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #72030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #72070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #72110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #72150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #72190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #72230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #72270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #72310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #72350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #72390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #72430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #72470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #72510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #72550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #72590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #72630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #72670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #72710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #72750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #72790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #72830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #72870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #72910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #72950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #72990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #73030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #73070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #73110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #73150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #73190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #73230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #73270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #73310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #73350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #73390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #73430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #73470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #73510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #73550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #73590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #73630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #73670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #73710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #73750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #73790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #73830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #73870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #73910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #73950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #73990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #74030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #74070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #74110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #74150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #74190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #74230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #74270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #74310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #74350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};
         #74390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd10, 4'd 4};
         #74430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd10, 4'd 4};
         #74470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd14, 4'd 4};
         #74510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd14, 4'd 4};
         #74550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 2, 4'd 4};
         #74590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 2, 4'd 4};
         #74630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 6, 4'd 4};
         #74670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 6, 4'd 4};
         #74710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd10, 4'd 4};
         #74750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd10, 4'd 4};
         #74790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd14, 4'd 4};
         #74830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd14, 4'd 4};
         #74870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 2, 4'd 4};
         #74910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 2, 4'd 4};
         #74950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 6, 4'd 4};
         #74990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 6, 4'd 4};

         #75000 {hsync, vsync, red, green, blue} <= {2'bxx, 4'd x, 4'd x, 4'd x};

         #16702070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16730230 {hsync, vsync, red, green, blue} <= {2'b01, 4'd 0, 4'd 0, 4'd 0};
         #16734070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16762230 {hsync, vsync, red, green, blue} <= {2'b01, 4'd 0, 4'd 0, 4'd 0};
         #16766070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16794230 {hsync, vsync, red, green, blue} <= {2'b01, 4'd 0, 4'd 0, 4'd 0};
         #16798070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16800030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16800070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16800110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16800150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16800190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16800230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16800270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16800310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16800350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16800390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16800430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16800470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16800510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16800550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16800590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16800630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16800670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16800710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16800750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16800790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16800830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16800870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16800910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16800950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16800990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16801030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16801070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16801110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16801150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16801190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16801230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16801270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16801310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16801350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16801390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16801430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16801470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16801510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16801550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16801590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16801630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16801670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16801710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16801750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16801790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16801830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16801870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16801910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16801950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16801990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16802030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16802070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16802110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16802150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16802190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16802230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16802270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16802310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16802350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16802390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16802430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16802470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16802510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16802550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16802590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16802630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16802670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16802710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16802750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16802790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16802830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16802870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16802910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16802950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16802990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16803030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16803070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16803110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16803150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16803190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16803230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16803270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16803310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16803350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16803390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16803430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16803470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16803510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16803550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16803590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16803630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16803670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16803710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16803750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16803790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16803830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16803870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16803910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16803950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16803990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16804030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16804070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16804110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16804150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16804190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16804230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16804270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16804310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16804350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16804390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16804430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16804470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16804510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16804550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16804590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16804630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16804670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16804710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16804750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16804790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16804830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16804870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16804910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16804950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16804990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16805030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16805070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16805110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16805150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16805190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16805230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16805270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16805310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16805350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16805390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16805430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16805470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16805510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16805550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16805590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16805630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16805670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16805710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16805750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16805790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16805830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16805870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16805910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16805950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16805990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16806030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16806070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16806110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16806150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16806190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16806230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16806270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16806310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16806350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16806390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16806430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16806470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16806510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16806550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16806590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16806630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16806670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16806710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16806750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16806790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16806830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16806870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16806910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16806950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16806990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16807030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16807070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16807110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16807150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16807190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16807230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16807270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16807310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16807350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16807390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16807430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16807470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16807510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16807550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16807590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16807630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16807670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16807710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16807750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16807790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16807830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16807870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16807910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16807950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16807990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16808030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16808070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16808110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16808150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16808190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16808230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16808270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16808310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16808350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16808390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16808430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16808470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16808510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16808550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16808590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16808630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16808670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16808710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16808750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16808790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16808830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16808870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16808910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16808950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16808990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16809030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16809070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16809110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16809150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16809190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16809230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16809270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16809310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16809350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16809390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16809430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16809470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16809510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16809550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16809590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16809630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16809670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16809710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16809750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16809790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16809830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16809870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16809910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16809950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16809990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16810030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16810070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16810110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16810150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16810190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16810230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16810270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16810310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16810350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16810390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16810430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16810470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16810510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16810550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16810590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16810630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16810670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16810710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16810750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16810790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16810830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16810870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16810910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16810950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16810990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16811030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16811070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16811110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16811150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16811190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16811230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16811270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16811310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16811350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16811390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16811430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16811470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16811510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16811550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16811590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16811630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16811670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16811710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16811750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16811790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16811830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16811870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16811910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16811950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16811990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16812030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16812070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16812110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16812150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16812190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16812230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16812270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16812310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16812350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16812390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16812430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16812470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16812510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16812550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16812590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16812630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16812670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16812710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16812750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16812790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16812830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16812870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16812910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16812950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16812990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16813030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16813070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16813110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16813150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16813190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16813230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16813270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16813310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16813350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16813390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16813430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16813470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16813510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16813550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16813590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16813630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16813670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16813710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16813750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16813790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16813830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16813870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16813910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16813950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16813990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16814030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16814070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16814110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16814150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16814190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16814230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16814270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16814310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16814350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16814390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16814430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16814470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16814510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16814550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16814590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16814630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16814670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16814710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16814750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16814790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16814830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16814870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16814910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16814950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16814990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16815030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16815070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16815110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16815150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16815190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16815230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16815270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16815310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16815350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16815390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16815430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16815470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16815510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16815550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16815590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16815630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16815670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16815710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16815750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16815790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16815830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16815870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16815910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16815950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16815990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16816030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16816070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16816110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16816150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16816190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16816230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16816270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16816310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16816350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16816390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16816430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16816470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16816510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16816550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16816590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16816630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16816670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16816710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16816750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16816790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16816830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16816870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16816910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16816950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16816990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16817030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16817070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16817110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16817150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16817190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16817230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16817270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16817310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16817350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16817390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16817430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16817470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16817510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16817550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16817590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16817630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16817670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16817710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16817750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16817790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16817830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16817870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16817910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16817950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16817990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16818030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16818070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16818110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16818150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16818190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16818230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16818270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16818310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16818350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16818390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16818430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16818470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16818510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16818550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16818590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16818630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16818670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16818710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16818750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16818790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16818830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16818870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16818910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16818950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16818990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16819030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16819070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16819110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16819150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16819190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16819230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16819270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16819310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16819350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16819390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16819430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16819470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16819510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16819550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16819590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16819630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16819670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16819710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16819750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16819790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16819830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16819870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16819910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16819950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16819990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16820030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16820070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16820110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16820150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16820190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16820230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16820270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16820310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16820350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16820390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16820430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16820470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16820510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16820550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16820590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16820630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16820670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16820710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16820750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16820790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16820830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16820870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16820910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16820950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16820990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16821030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16821070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16821110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16821150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16821190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16821230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16821270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16821310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16821350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16821390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16821430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16821470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16821510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16821550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16821590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16821630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16821670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16821710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16821750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16821790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16821830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16821870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16821910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16821950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16821990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16822030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16822070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16822110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16822150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16822190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16822230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16822270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16822310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16822350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16822390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16822430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16822470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16822510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16822550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16822590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16822630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16822670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16822710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16822750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16822790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16822830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16822870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16822910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16822950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16822990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16823030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16823070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16823110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16823150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16823190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16823230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16823270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16823310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16823350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16823390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16823430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16823470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16823510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16823550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16823590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16823630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16823670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16823710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16823750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16823790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16823830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16823870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16823910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16823950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16823990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16824030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16824070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16824110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16824150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16824190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16824230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16824270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16824310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16824350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16824390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16824430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16824470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16824510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16824550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16824590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16824630 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16824670 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16824710 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16824750 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16824790 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16824830 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16824870 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16824910 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16824950 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16824990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 1, 4'd 0, 4'd 0};
         #16825030 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 2, 4'd 4, 4'd 0};
         #16825070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 3, 4'd 4, 4'd 0};
         #16825110 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 4, 4'd 8, 4'd 0};
         #16825150 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 5, 4'd 8, 4'd 0};
         #16825190 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 6, 4'd12, 4'd 0};
         #16825230 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 7, 4'd12, 4'd 0};
         #16825270 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 8, 4'd 0, 4'd 0};
         #16825310 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 9, 4'd 0, 4'd 0};
         #16825350 {hsync, vsync, red, green, blue} <= {2'b11, 4'd10, 4'd 4, 4'd 0};
         #16825390 {hsync, vsync, red, green, blue} <= {2'b11, 4'd11, 4'd 4, 4'd 0};
         #16825430 {hsync, vsync, red, green, blue} <= {2'b11, 4'd12, 4'd 8, 4'd 0};
         #16825470 {hsync, vsync, red, green, blue} <= {2'b11, 4'd13, 4'd 8, 4'd 0};
         #16825510 {hsync, vsync, red, green, blue} <= {2'b11, 4'd14, 4'd12, 4'd 0};
         #16825550 {hsync, vsync, red, green, blue} <= {2'b11, 4'd15, 4'd12, 4'd 0};
         #16825590 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16826230 {hsync, vsync, red, green, blue} <= {2'b01, 4'd 0, 4'd 0, 4'd 0};
         #16830070 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 0, 4'd 0};
         #16831990 {hsync, vsync, red, green, blue} <= {2'b11, 4'd 0, 4'd 1, 4'd 2};
      join
   end
endmodule